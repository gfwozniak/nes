package Games;

typedef enum logic [3:0] {MARIO, DONKEY_KONG, NES_TEST} game_name;

endpackage : Games